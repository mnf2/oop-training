`ifndef TOP
`define TOP

module top();
    initial begin

        // Add your code here.

        // Finish the test.
        $finish();
    end
endmodule

`endif // TOP
